----------------------------------------------------------------------------------
-- Company: USAFA
-- Engineer: C3C Combs
-- 
-- Create Date:    10:33:47 07/07/2012 
-- Design Name: 
-- Module Name:    MooreElevatorController_Silva - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: This is the component code for a Mealy Elevator.  The inputs directly affect the outputs.
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MealyElevatorController_Shell is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           stop : in  STD_LOGIC;
           up_down : in  STD_LOGIC;
           floorOne : out  STD_LOGIC_VECTOR (3 downto 0);
			  floorTen : out STD_LOGIC_VECTOR (3 downto 0);
			  nextfloor : out std_logic_vector (3 downto 0));
end MealyElevatorController_Shell;

architecture Behavioral of MealyElevatorController_Shell is

type floor_state_type is (floor1, floor2, floor3, floor4, floor5, floor6, floor7, floor8, floor9, floor10, floor11, floor12, floor13, floor14, floor15, floor16, floor17, floor18, floor19, floor20, floor21, floor22, floor23);

signal floor_state : floor_state_type;

begin

---------------------------------------------------------
--Code your Mealy machine next-state process below
--Question: Will it be different from your Moore Machine?
---------------------------------------------------------
floor_state_machine: process(clk)
begin
	--clk'event and clk='1' is VHDL-speak for a rising edge
	if clk'event and clk='1' then
		--reset is active high and will return the elevator to floor1
		--Question: is reset synchronous or asynchronous?
		if reset='1' then
			floor_state <= floor1;
		--now we will code our next-state logic
		else
			case floor_state is
				--when our current state is floor1
				when floor1 =>
					--if up_down is set to "go up" and stop is set to 
					--"don't stop" which floor do we want to go to?
					if (up_down='1' and stop='0') then 
						--floor2 right?? This makes sense!
						floor_state <= floor2;
					--otherwise we're going to stay at floor1
					else
						floor_state <= floor1;
					end if;
				--when our current state is floor2
				when floor2 => 
					--if up_down is set to "go up" and stop is set to 
					--"don't stop" which floor do we want to go to?
					if (up_down='1' and stop='0') then 
						floor_state <= floor3; 			
					--if up_down is set to "go down" and stop is set to 
					--"don't stop" which floor do we want to go to?
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor1;
					--otherwise we're going to stay at floor2
					else
						floor_state <= floor2;
					end if;
				
--COMPLETE THE NEXT STATE LOGIC ASSIGNMENTS FOR FLOORS 3 AND 4
				when floor3 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor4;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor2;	
					else
						floor_state <= floor3;	
					end if;
				when floor4 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor5;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor3;	
					else
						floor_state <= floor4;	
					end if;
				when floor5 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor6;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor4;	
					else
						floor_state <= floor5;	
					end if;
				when floor6 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor7;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor5;	
					else
						floor_state <= floor6;	
					end if;
				when floor7 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor8;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor6;	
					else
						floor_state <= floor7;	
					end if;
				when floor8 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor9;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor7;	
					else
						floor_state <= floor8;	
					end if;
				when floor9 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor10;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor8;	
					else
						floor_state <= floor9;	
					end if;
				when floor10 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor11;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor9;	
					else
						floor_state <= floor10;	
					end if;
				when floor11 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor12;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor10;	
					else
						floor_state <= floor11;	
					end if;
				when floor12 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor13;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor11;	
					else
						floor_state <= floor12;	
					end if;
				when floor13 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor14;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor12;	
					else
						floor_state <= floor13;	
					end if;
				when floor14 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor15;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor13;	
					else
						floor_state <= floor14;	
					end if;
				when floor15 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor15;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor14;	
					else
						floor_state <= floor15;	
					end if;	
				--This line accounts for phantom states
				when others =>
					floor_state <= floor1;
			end case;
		end if;
	end if;
end process;

-----------------------------------------------------------
--Code your Ouput Logic for your Mealy machine below
--Remember, now you have 2 outputs (floor and nextfloor)
-----------------------------------------------------------
floorOne <= "0001" when (floor_state = floor1) else
			"0010" when (floor_state = floor2) else
			"0011" when (floor_state = floor3) else
			"0100" when (floor_state = floor4) else
			"0101" when (floor_state = floor5) else
			"0110" when (floor_state = floor6) else
			"0111" when (floor_state = floor7) else
			"1000" when (floor_state = floor8) else
			"1001" when (floor_state = floor9) else
			"0000" when (floor_state = floor10) else
			"0001" when (floor_state = floor11) else
			"0010" when (floor_state = floor12) else
			"0011" when (floor_state = floor13) else
			"0100" when (floor_state = floor14) else
			"0101" when (floor_state = floor15) else
			"0001";
floorTen <= "0000" when (floor_state = floor1) else
			"0000" when (floor_state = floor2) else
			"0000" when (floor_state = floor3) else
			"0000" when (floor_state = floor4) else
			"0000" when (floor_state = floor5) else
			"0000" when (floor_state = floor6) else
			"0000" when (floor_state = floor7) else
			"0000" when (floor_state = floor8) else
			"0000" when (floor_state = floor9) else
			"0001" when (floor_state = floor10) else
			"0001" when (floor_state = floor11) else
			"0001" when (floor_state = floor12) else
			"0001" when (floor_state = floor13) else
			"0001" when (floor_state = floor14) else
			"0001" when (floor_state = floor15) else
			"0000";
nextfloor <= "0001" when ((floor_state = floor1 and up_down = '0') or reset = '1') else
			"0010" when ((floor_state = floor2 and stop = '1') or (floor_state = floor1 and up_down = '1' and stop = '0') or (floor_state = floor3 and up_down = '0' and stop = '0')) else
			"0011" when ((floor_state = floor3 and stop = '1') or (floor_state = floor2 and up_down = '1' and stop = '0') or (floor_state = floor4 and up_down = '0' and stop = '0')) else
			"0100" when ((floor_state = floor4 and stop = '1') or (floor_state = floor3 and up_down = '1' and stop = '0') or (floor_state = floor5 and up_down = '0' and stop = '0')) else
			"0101" when ((floor_state = floor5 and stop = '1') or (floor_state = floor4 and up_down = '1' and stop = '0') or (floor_state = floor6 and up_down = '0' and stop = '0')) else
			"0110" when ((floor_state = floor6 and stop = '1') or (floor_state = floor5 and up_down = '1' and stop = '0') or (floor_state = floor7 and up_down = '0' and stop = '0')) else
			"0111" when ((floor_state = floor7 and stop = '1') or (floor_state = floor6 and up_down = '1' and stop = '0') or (floor_state = floor8 and up_down = '0' and stop = '0')) else
			"1000" when ((floor_state = floor8 and stop = '1') or (floor_state = floor7 and up_down = '1' and stop = '0') or (floor_state = floor9 and up_down = '0' and stop = '0')) else
			"1001" when ((floor_state = floor9 and stop = '1') or (floor_state = floor8 and up_down = '1' and stop = '0') or (floor_state = floor10 and up_down = '0' and stop = '0')) else
			"1010" when ((floor_state = floor10 and stop = '1') or (floor_state = floor9 and up_down = '1' and stop = '0') or (floor_state = floor11 and up_down = '0' and stop = '0')) else
			"1011" when ((floor_state = floor11 and stop = '1') or (floor_state = floor10 and up_down = '1' and stop = '0') or (floor_state = floor12 and up_down = '0' and stop = '0')) else
			"1100" when ((floor_state = floor12 and stop = '1') or (floor_state = floor11 and up_down = '1' and stop = '0') or (floor_state = floor13 and up_down = '0' and stop = '0')) else
			"1101" when ((floor_state = floor13 and stop = '1') or (floor_state = floor12 and up_down = '1' and stop = '0') or (floor_state = floor14 and up_down = '0' and stop = '0')) else
			"1110" when ((floor_state = floor14 and stop = '1') or (floor_state = floor13 and up_down = '1' and stop = '0') or (floor_state = floor15 and up_down = '0' and stop = '0')) else
			"1111" when ((floor_state = floor15 and stop = '1') or (floor_state = floor14 and up_down = '1' and stop = '0')) else
			"0001";	

end Behavioral;

