----------------------------------------------------------------------------------
-- Company: USAFA
-- Engineer: C3C Combs
-- 
-- Create Date:    	10:33:47 07/07/2012 
-- Design Name:		CE3
-- Module Name:    	MooreElevatorController_Shell - Behavioral 
-- Description: 		Component code for a Moore Elevator machine.
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MooreElevatorController_Shell is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           stop : in  STD_LOGIC;
           up_down : in  STD_LOGIC;
           floorOne : out  STD_LOGIC_VECTOR (3 downto 0);
			  floorTen : out STD_LOGIC_VECTOR (3 downto 0);
			  LEDO : out STD_LOGIC_VECTOR (7 downto 0));
end MooreElevatorController_Shell;

architecture Behavioral of MooreElevatorController_Shell is

--Below you create a new variable type! You also define what values that 
--variable type can take on. Now you can assign a signal as 
--"floor_state_type" the same way you'd assign a signal as std_logic 
type floor_state_type is (floor1, floor2, floor3, floor4, floor5, floor6, floor7, floor8, floor9, floor10, floor11, floor12, floor13, floor14, floor15, floor16, floor17, floor18, floor19, floor20, floor21, floor22, floor23);

--Here you create a variable "floor_state" that can take on the values
--defined above. Neat-o!
signal floor_state : floor_state_type;

begin
---------------------------------------------
--Below you will code your next-state process
---------------------------------------------

--This line will set up a process that is sensitive to the clock
floor_state_machine: process(clk)
begin
	--clk'event and clk='1' is VHDL-speak for a rising edge
	if clk'event and clk='1' then
		--reset is active high and will return the elevator to floor1
		--Question: is reset synchronous or asynchronous?
		if reset='1' then
			floor_state <= floor1;
		--now we will code our next-state logic
		else
			case floor_state is
				--when our current state is floor1
				when floor1 =>
					--if up_down is set to "go up" and stop is set to 
					--"don't stop" which floor do we want to go to?
					if (up_down='1' and stop='0') then 
						--floor2 right?? This makes sense!
						floor_state <= floor2;
					--otherwise we're going to stay at floor1
					else
						floor_state <= floor1;
					end if;
				--when our current state is floor2
				when floor2 => 
					--if up_down is set to "go up" and stop is set to 
					--"don't stop" which floor do we want to go to?
					if (up_down='1' and stop='0') then 
						floor_state <= floor3; 			
					--if up_down is set to "go down" and stop is set to 
					--"don't stop" which floor do we want to go to?
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor1;
					--otherwise we're going to stay at floor2
					else
						floor_state <= floor2;
					end if;
				
--COMPLETE THE NEXT STATE LOGIC ASSIGNMENTS FOR FLOORS 3 AND 4
				when floor3 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor4;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor2;	
					else
						floor_state <= floor3;	
					end if;
				when floor4 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor5;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor3;	
					else
						floor_state <= floor4;	
					end if;
				when floor5 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor6;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor4;	
					else
						floor_state <= floor5;	
					end if;
				when floor6 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor7;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor5;	
					else
						floor_state <= floor6;	
					end if;
				when floor7 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor8;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor6;	
					else
						floor_state <= floor7;	
					end if;
				when floor8 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor9;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor7;	
					else
						floor_state <= floor8;	
					end if;
				when floor9 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor10;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor8;	
					else
						floor_state <= floor9;	
					end if;
				when floor10 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor11;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor9;	
					else
						floor_state <= floor10;	
					end if;
				when floor11 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor12;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor10;	
					else
						floor_state <= floor11;	
					end if;
				when floor12 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor13;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor11;	
					else
						floor_state <= floor12;	
					end if;
				when floor13 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor14;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor12;	
					else
						floor_state <= floor13;	
					end if;
				when floor14 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor15;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor13;	
					else
						floor_state <= floor14;	
					end if;
				when floor15 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor16;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor14;	
					else
						floor_state <= floor15;	
					end if;
				when floor16 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor17;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor15;	
					else
						floor_state <= floor16;	
					end if;
				when floor17 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor18;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor16;	
					else
						floor_state <= floor17;	
					end if;
				when floor18 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor19;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor17;	
					else
						floor_state <= floor18;	
					end if;
				when floor19 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor20;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor18;	
					else
						floor_state <= floor19;	
					end if;
				when floor20 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor21;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor19;	
					else
						floor_state <= floor20;	
					end if;
				when floor21 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor22;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor20;	
					else
						floor_state <= floor21;	
					end if;
				when floor22 =>
					if (up_down='1' and stop='0') then 
						floor_state <= floor23;
					elsif (up_down='0' and stop='0') then 
						floor_state <= floor21;	
					else
						floor_state <= floor22;	
					end if;
				when floor23 =>
					if (up_down='0' and stop='0') then 
						floor_state <= floor22;	
					else
						floor_state <= floor23;	
					end if;
				
				--This line accounts for phantom states
				when others =>
					floor_state <= floor1;
			end case;
		end if;
	end if;
end process;
-- Here you define your output logic. Finish the statements below
floorOne <= "0001" when (floor_state = floor1) else
			"0010" when (floor_state = floor2) else
			"0011" when (floor_state = floor3) else
			"0100" when (floor_state = floor4) else
			"0101" when (floor_state = floor5) else
			"0110" when (floor_state = floor6) else
			"0111" when (floor_state = floor7) else
			"1000" when (floor_state = floor8) else
			"1001" when (floor_state = floor9) else
			"0000" when (floor_state = floor10) else
			"0001" when (floor_state = floor11) else
			"0010" when (floor_state = floor12) else
			"0011" when (floor_state = floor13) else
			"0100" when (floor_state = floor14) else
			"0101" when (floor_state = floor15) else
			"0110" when (floor_state = floor16) else
			"0111" when (floor_state = floor17) else
			"1000" when (floor_state = floor18) else
			"1001" when (floor_state = floor19) else
			"0000" when (floor_state = floor20) else
			"0001" when (floor_state = floor21) else
			"0010" when (floor_state = floor22) else
			"0011" when (floor_state = floor23) else
			"0010";
floorTen <= "0000" when (floor_state = floor1) else
			"0000" when (floor_state = floor2) else
			"0000" when (floor_state = floor3) else
			"0000" when (floor_state = floor4) else
			"0000" when (floor_state = floor5) else
			"0000" when (floor_state = floor6) else
			"0000" when (floor_state = floor7) else
			"0000" when (floor_state = floor8) else
			"0000" when (floor_state = floor9) else
			"0001" when (floor_state = floor10) else
			"0001" when (floor_state = floor11) else
			"0001" when (floor_state = floor12) else
			"0001" when (floor_state = floor13) else
			"0001" when (floor_state = floor14) else
			"0001" when (floor_state = floor15) else
			"0001" when (floor_state = floor16) else
			"0001" when (floor_state = floor17) else
			"0001" when (floor_state = floor18) else
			"0001" when (floor_state = floor19) else
			"0010" when (floor_state = floor20) else
			"0010" when (floor_state = floor21) else
			"0010" when (floor_state = floor22) else
			"0010" when (floor_state = floor23) else
			"0000";
LEDO <= "00000001" when (floor_state = floor1) else
         "00000010" when (floor_state = floor2) else
			"00000100" when (floor_state = floor3) else
			"00001000" when (floor_state = floor4) else
			"00010000" when (floor_state = floor5) else
			"00100000" when (floor_state = floor6) else
			"01000000" when (floor_state = floor7) else
			"10000000" when (floor_state = floor8) else
			"00000001" when (floor_state = floor9) else
			"00000010" when (floor_state = floor10) else
			"00000100" when (floor_state = floor11) else
			"00001000" when (floor_state = floor12) else
			"00010000" when (floor_state = floor13) else
			"00100000" when (floor_state = floor14) else
			"01000000" when (floor_state = floor15) else
			"10000000" when (floor_state = floor16) else
			"00000001" when (floor_state = floor17) else
			"00000010" when (floor_state = floor18) else
			"00000100" when (floor_state = floor19) else
			"00001000" when (floor_state = floor20) else
			"00010000" when (floor_state = floor21) else
			"00100000" when (floor_state = floor22) else
			"01000000" when (floor_state = floor23) else
			"00000001";
end Behavioral;

